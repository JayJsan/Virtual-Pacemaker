// nios2_system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module nios2_system (
		input  wire        clk_clk,                               //                            clk.clk
		input  wire [2:0]  keys_external_connection_export,       //       keys_external_connection.export
		output wire        lcd_external_RS,                       //                   lcd_external.RS
		output wire        lcd_external_RW,                       //                               .RW
		inout  wire [7:0]  lcd_external_data,                     //                               .data
		output wire        lcd_external_E,                        //                               .E
		output wire [8:0]  leds_green_external_connection_export, // leds_green_external_connection.export
		output wire [17:0] leds_red_external_connection_export,   //   leds_red_external_connection.export
		input  wire        reset_reset_n,                         //                          reset.reset_n
		output wire        sdram_pll_sdram_clk_clk,               //            sdram_pll_sdram_clk.clk
		output wire [11:0] sdram_wire_addr,                       //                     sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                         //                               .ba
		output wire        sdram_wire_cas_n,                      //                               .cas_n
		output wire        sdram_wire_cke,                        //                               .cke
		output wire        sdram_wire_cs_n,                       //                               .cs_n
		inout  wire [15:0] sdram_wire_dq,                         //                               .dq
		output wire [1:0]  sdram_wire_dqm,                        //                               .dqm
		output wire        sdram_wire_ras_n,                      //                               .ras_n
		output wire        sdram_wire_we_n,                       //                               .we_n
		input  wire [17:0] switches_external_connection_export,   //   switches_external_connection.export
		input  wire        uart_external_connection_rxd,          //       uart_external_connection.rxd
		output wire        uart_external_connection_txd           //                               .txd
	);

	wire         sdram_pll_sys_clk_clk;                                     // sdram_pll:sys_clk_clk -> [cpu:clk, irq_mapper:clk, jtag_uart:clk, keys:clk, lcd:clk, leds_green:clk, leds_red:clk, mm_interconnect_0:sdram_pll_sys_clk_clk, onchip_mem:clk, rst_controller:clk, sdram:clk, switches:clk, timer_0:clk, timer_1:clk, uart:clk]
	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [24:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                             // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [24:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                      // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [7:0] mm_interconnect_0_lcd_control_slave_readdata;              // lcd:readdata -> mm_interconnect_0:lcd_control_slave_readdata
	wire   [1:0] mm_interconnect_0_lcd_control_slave_address;               // mm_interconnect_0:lcd_control_slave_address -> lcd:address
	wire         mm_interconnect_0_lcd_control_slave_read;                  // mm_interconnect_0:lcd_control_slave_read -> lcd:read
	wire         mm_interconnect_0_lcd_control_slave_begintransfer;         // mm_interconnect_0:lcd_control_slave_begintransfer -> lcd:begintransfer
	wire         mm_interconnect_0_lcd_control_slave_write;                 // mm_interconnect_0:lcd_control_slave_write -> lcd:write
	wire   [7:0] mm_interconnect_0_lcd_control_slave_writedata;             // mm_interconnect_0:lcd_control_slave_writedata -> lcd:writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_mem_s1_chipselect;                // mm_interconnect_0:onchip_mem_s1_chipselect -> onchip_mem:chipselect
	wire  [15:0] mm_interconnect_0_onchip_mem_s1_readdata;                  // onchip_mem:readdata -> mm_interconnect_0:onchip_mem_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_mem_s1_address;                   // mm_interconnect_0:onchip_mem_s1_address -> onchip_mem:address
	wire   [1:0] mm_interconnect_0_onchip_mem_s1_byteenable;                // mm_interconnect_0:onchip_mem_s1_byteenable -> onchip_mem:byteenable
	wire         mm_interconnect_0_onchip_mem_s1_write;                     // mm_interconnect_0:onchip_mem_s1_write -> onchip_mem:write
	wire  [15:0] mm_interconnect_0_onchip_mem_s1_writedata;                 // mm_interconnect_0:onchip_mem_s1_writedata -> onchip_mem:writedata
	wire         mm_interconnect_0_onchip_mem_s1_clken;                     // mm_interconnect_0:onchip_mem_s1_clken -> onchip_mem:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_uart_s1_chipselect;                      // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                        // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                         // mm_interconnect_0:uart_s1_address -> uart:address
	wire         mm_interconnect_0_uart_s1_read;                            // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;                   // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                           // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                       // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                   // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                     // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                      // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                        // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                    // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_timer_1_s1_chipselect;                   // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                     // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                      // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                        // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                    // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire         mm_interconnect_0_keys_s1_chipselect;                      // mm_interconnect_0:keys_s1_chipselect -> keys:chipselect
	wire  [31:0] mm_interconnect_0_keys_s1_readdata;                        // keys:readdata -> mm_interconnect_0:keys_s1_readdata
	wire   [1:0] mm_interconnect_0_keys_s1_address;                         // mm_interconnect_0:keys_s1_address -> keys:address
	wire         mm_interconnect_0_keys_s1_write;                           // mm_interconnect_0:keys_s1_write -> keys:write_n
	wire  [31:0] mm_interconnect_0_keys_s1_writedata;                       // mm_interconnect_0:keys_s1_writedata -> keys:writedata
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                    // switches:readdata -> mm_interconnect_0:switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                     // mm_interconnect_0:switches_s1_address -> switches:address
	wire         mm_interconnect_0_leds_red_s1_chipselect;                  // mm_interconnect_0:leds_red_s1_chipselect -> leds_red:chipselect
	wire  [31:0] mm_interconnect_0_leds_red_s1_readdata;                    // leds_red:readdata -> mm_interconnect_0:leds_red_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_red_s1_address;                     // mm_interconnect_0:leds_red_s1_address -> leds_red:address
	wire         mm_interconnect_0_leds_red_s1_write;                       // mm_interconnect_0:leds_red_s1_write -> leds_red:write_n
	wire  [31:0] mm_interconnect_0_leds_red_s1_writedata;                   // mm_interconnect_0:leds_red_s1_writedata -> leds_red:writedata
	wire         mm_interconnect_0_leds_green_s1_chipselect;                // mm_interconnect_0:leds_green_s1_chipselect -> leds_green:chipselect
	wire  [31:0] mm_interconnect_0_leds_green_s1_readdata;                  // leds_green:readdata -> mm_interconnect_0:leds_green_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_green_s1_address;                   // mm_interconnect_0:leds_green_s1_address -> leds_green:address
	wire         mm_interconnect_0_leds_green_s1_write;                     // mm_interconnect_0:leds_green_s1_write -> leds_green:write_n
	wire  [31:0] mm_interconnect_0_leds_green_s1_writedata;                 // mm_interconnect_0:leds_green_s1_writedata -> leds_green:writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // timer_1:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // timer_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // keys:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                  // uart:irq -> irq_mapper:receiver4_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [cpu:reset_n, irq_mapper:reset, jtag_uart:rst_n, keys:reset_n, lcd:reset_n, leds_green:reset_n, leds_red:reset_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchip_mem:reset, rst_translator:in_reset, sdram:reset_n, switches:reset_n, timer_0:reset_n, timer_1:reset_n, uart:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, onchip_mem:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> sdram_pll:ref_reset_reset

	nios2_system_cpu cpu (
		.clk                                 (sdram_pll_sys_clk_clk),                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	nios2_system_jtag_uart jtag_uart (
		.clk            (sdram_pll_sys_clk_clk),                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	nios2_system_keys keys (
		.clk        (sdram_pll_sys_clk_clk),                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_keys_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keys_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keys_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keys_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keys_s1_readdata),   //                    .readdata
		.in_port    (keys_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver3_irq)              //                 irq.irq
	);

	nios2_system_lcd lcd (
		.reset_n       (~rst_controller_reset_out_reset),                   //         reset.reset_n
		.clk           (sdram_pll_sys_clk_clk),                             //           clk.clk
		.begintransfer (mm_interconnect_0_lcd_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_0_lcd_control_slave_read),          //              .read
		.write         (mm_interconnect_0_lcd_control_slave_write),         //              .write
		.readdata      (mm_interconnect_0_lcd_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_0_lcd_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_0_lcd_control_slave_address),       //              .address
		.LCD_RS        (lcd_external_RS),                                   //      external.export
		.LCD_RW        (lcd_external_RW),                                   //              .export
		.LCD_data      (lcd_external_data),                                 //              .export
		.LCD_E         (lcd_external_E)                                     //              .export
	);

	nios2_system_leds_green leds_green (
		.clk        (sdram_pll_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_leds_green_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_green_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_green_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_green_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_green_s1_readdata),   //                    .readdata
		.out_port   (leds_green_external_connection_export)       // external_connection.export
	);

	nios2_system_leds_red leds_red (
		.clk        (sdram_pll_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_leds_red_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_red_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_red_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_red_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_red_s1_readdata),   //                    .readdata
		.out_port   (leds_red_external_connection_export)       // external_connection.export
	);

	nios2_system_onchip_mem onchip_mem (
		.clk        (sdram_pll_sys_clk_clk),                      //   clk1.clk
		.address    (mm_interconnect_0_onchip_mem_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_mem_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_mem_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_mem_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_mem_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_mem_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_mem_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	nios2_system_sdram sdram (
		.clk            (sdram_pll_sys_clk_clk),                    //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	nios2_system_sdram_pll sdram_pll (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (rst_controller_001_reset_out_reset), //    ref_reset.reset
		.sys_clk_clk        (sdram_pll_sys_clk_clk),              //      sys_clk.clk
		.sdram_clk_clk      (sdram_pll_sdram_clk_clk),            //    sdram_clk.clk
		.reset_source_reset ()                                    // reset_source.reset
	);

	nios2_system_switches switches (
		.clk      (sdram_pll_sys_clk_clk),                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_external_connection_export)     // external_connection.export
	);

	nios2_system_timer_0 timer_0 (
		.clk        (sdram_pll_sys_clk_clk),                   //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                 //   irq.irq
	);

	nios2_system_timer_0 timer_1 (
		.clk        (sdram_pll_sys_clk_clk),                   //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	nios2_system_uart uart (
		.clk           (sdram_pll_sys_clk_clk),                   //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.endofpacket   (),                                        //                    .endofpacket
		.rxd           (uart_external_connection_rxd),            // external_connection.export
		.txd           (uart_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver4_irq)                 //                 irq.irq
	);

	nios2_system_mm_interconnect_0 mm_interconnect_0 (
		.sdram_pll_sys_clk_clk                   (sdram_pll_sys_clk_clk),                                     //               sdram_pll_sys_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                            // cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                 (cpu_data_master_address),                                   //                 cpu_data_master.address
		.cpu_data_master_waitrequest             (cpu_data_master_waitrequest),                               //                                .waitrequest
		.cpu_data_master_byteenable              (cpu_data_master_byteenable),                                //                                .byteenable
		.cpu_data_master_read                    (cpu_data_master_read),                                      //                                .read
		.cpu_data_master_readdata                (cpu_data_master_readdata),                                  //                                .readdata
		.cpu_data_master_readdatavalid           (cpu_data_master_readdatavalid),                             //                                .readdatavalid
		.cpu_data_master_write                   (cpu_data_master_write),                                     //                                .write
		.cpu_data_master_writedata               (cpu_data_master_writedata),                                 //                                .writedata
		.cpu_data_master_debugaccess             (cpu_data_master_debugaccess),                               //                                .debugaccess
		.cpu_instruction_master_address          (cpu_instruction_master_address),                            //          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest      (cpu_instruction_master_waitrequest),                        //                                .waitrequest
		.cpu_instruction_master_read             (cpu_instruction_master_read),                               //                                .read
		.cpu_instruction_master_readdata         (cpu_instruction_master_readdata),                           //                                .readdata
		.cpu_instruction_master_readdatavalid    (cpu_instruction_master_readdatavalid),                      //                                .readdatavalid
		.cpu_debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),             //             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                .write
		.cpu_debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                .read
		.cpu_debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                .readdata
		.cpu_debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                .writedata
		.cpu_debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                .byteenable
		.cpu_debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                .waitrequest
		.cpu_debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                .debugaccess
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                .chipselect
		.keys_s1_address                         (mm_interconnect_0_keys_s1_address),                         //                         keys_s1.address
		.keys_s1_write                           (mm_interconnect_0_keys_s1_write),                           //                                .write
		.keys_s1_readdata                        (mm_interconnect_0_keys_s1_readdata),                        //                                .readdata
		.keys_s1_writedata                       (mm_interconnect_0_keys_s1_writedata),                       //                                .writedata
		.keys_s1_chipselect                      (mm_interconnect_0_keys_s1_chipselect),                      //                                .chipselect
		.lcd_control_slave_address               (mm_interconnect_0_lcd_control_slave_address),               //               lcd_control_slave.address
		.lcd_control_slave_write                 (mm_interconnect_0_lcd_control_slave_write),                 //                                .write
		.lcd_control_slave_read                  (mm_interconnect_0_lcd_control_slave_read),                  //                                .read
		.lcd_control_slave_readdata              (mm_interconnect_0_lcd_control_slave_readdata),              //                                .readdata
		.lcd_control_slave_writedata             (mm_interconnect_0_lcd_control_slave_writedata),             //                                .writedata
		.lcd_control_slave_begintransfer         (mm_interconnect_0_lcd_control_slave_begintransfer),         //                                .begintransfer
		.leds_green_s1_address                   (mm_interconnect_0_leds_green_s1_address),                   //                   leds_green_s1.address
		.leds_green_s1_write                     (mm_interconnect_0_leds_green_s1_write),                     //                                .write
		.leds_green_s1_readdata                  (mm_interconnect_0_leds_green_s1_readdata),                  //                                .readdata
		.leds_green_s1_writedata                 (mm_interconnect_0_leds_green_s1_writedata),                 //                                .writedata
		.leds_green_s1_chipselect                (mm_interconnect_0_leds_green_s1_chipselect),                //                                .chipselect
		.leds_red_s1_address                     (mm_interconnect_0_leds_red_s1_address),                     //                     leds_red_s1.address
		.leds_red_s1_write                       (mm_interconnect_0_leds_red_s1_write),                       //                                .write
		.leds_red_s1_readdata                    (mm_interconnect_0_leds_red_s1_readdata),                    //                                .readdata
		.leds_red_s1_writedata                   (mm_interconnect_0_leds_red_s1_writedata),                   //                                .writedata
		.leds_red_s1_chipselect                  (mm_interconnect_0_leds_red_s1_chipselect),                  //                                .chipselect
		.onchip_mem_s1_address                   (mm_interconnect_0_onchip_mem_s1_address),                   //                   onchip_mem_s1.address
		.onchip_mem_s1_write                     (mm_interconnect_0_onchip_mem_s1_write),                     //                                .write
		.onchip_mem_s1_readdata                  (mm_interconnect_0_onchip_mem_s1_readdata),                  //                                .readdata
		.onchip_mem_s1_writedata                 (mm_interconnect_0_onchip_mem_s1_writedata),                 //                                .writedata
		.onchip_mem_s1_byteenable                (mm_interconnect_0_onchip_mem_s1_byteenable),                //                                .byteenable
		.onchip_mem_s1_chipselect                (mm_interconnect_0_onchip_mem_s1_chipselect),                //                                .chipselect
		.onchip_mem_s1_clken                     (mm_interconnect_0_onchip_mem_s1_clken),                     //                                .clken
		.sdram_s1_address                        (mm_interconnect_0_sdram_s1_address),                        //                        sdram_s1.address
		.sdram_s1_write                          (mm_interconnect_0_sdram_s1_write),                          //                                .write
		.sdram_s1_read                           (mm_interconnect_0_sdram_s1_read),                           //                                .read
		.sdram_s1_readdata                       (mm_interconnect_0_sdram_s1_readdata),                       //                                .readdata
		.sdram_s1_writedata                      (mm_interconnect_0_sdram_s1_writedata),                      //                                .writedata
		.sdram_s1_byteenable                     (mm_interconnect_0_sdram_s1_byteenable),                     //                                .byteenable
		.sdram_s1_readdatavalid                  (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                .readdatavalid
		.sdram_s1_waitrequest                    (mm_interconnect_0_sdram_s1_waitrequest),                    //                                .waitrequest
		.sdram_s1_chipselect                     (mm_interconnect_0_sdram_s1_chipselect),                     //                                .chipselect
		.switches_s1_address                     (mm_interconnect_0_switches_s1_address),                     //                     switches_s1.address
		.switches_s1_readdata                    (mm_interconnect_0_switches_s1_readdata),                    //                                .readdata
		.timer_0_s1_address                      (mm_interconnect_0_timer_0_s1_address),                      //                      timer_0_s1.address
		.timer_0_s1_write                        (mm_interconnect_0_timer_0_s1_write),                        //                                .write
		.timer_0_s1_readdata                     (mm_interconnect_0_timer_0_s1_readdata),                     //                                .readdata
		.timer_0_s1_writedata                    (mm_interconnect_0_timer_0_s1_writedata),                    //                                .writedata
		.timer_0_s1_chipselect                   (mm_interconnect_0_timer_0_s1_chipselect),                   //                                .chipselect
		.timer_1_s1_address                      (mm_interconnect_0_timer_1_s1_address),                      //                      timer_1_s1.address
		.timer_1_s1_write                        (mm_interconnect_0_timer_1_s1_write),                        //                                .write
		.timer_1_s1_readdata                     (mm_interconnect_0_timer_1_s1_readdata),                     //                                .readdata
		.timer_1_s1_writedata                    (mm_interconnect_0_timer_1_s1_writedata),                    //                                .writedata
		.timer_1_s1_chipselect                   (mm_interconnect_0_timer_1_s1_chipselect),                   //                                .chipselect
		.uart_s1_address                         (mm_interconnect_0_uart_s1_address),                         //                         uart_s1.address
		.uart_s1_write                           (mm_interconnect_0_uart_s1_write),                           //                                .write
		.uart_s1_read                            (mm_interconnect_0_uart_s1_read),                            //                                .read
		.uart_s1_readdata                        (mm_interconnect_0_uart_s1_readdata),                        //                                .readdata
		.uart_s1_writedata                       (mm_interconnect_0_uart_s1_writedata),                       //                                .writedata
		.uart_s1_begintransfer                   (mm_interconnect_0_uart_s1_begintransfer),                   //                                .begintransfer
		.uart_s1_chipselect                      (mm_interconnect_0_uart_s1_chipselect)                       //                                .chipselect
	);

	nios2_system_irq_mapper irq_mapper (
		.clk           (sdram_pll_sys_clk_clk),          //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (sdram_pll_sys_clk_clk),              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
